library ieee;
use ieee.std_logic_1164.all;

package Constants is
    
constant cHIGH  : std_logic := '1';
constant cHIGHN : std_logic := '0';
constant cLOW   : std_logic := '0';
constant cLOWN  : std_logic := '1';

constant cBYTELEN : integer := 8;
    
end package Constants;
