library ieee;
use ieee.std_logic_1164.all;

package Utilities is

function fNextpow2(a:in integer) return integer;

end package Utilities;

